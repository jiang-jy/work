/*
 *  TOPPERS/ASP Kernel
 *      Toyohashi Open Platform for Embedded Real-Time Systems/
 *      Advanced Standard Profile Kernel
 * 
 *  Copyright (C) 2015 by Ushio Laboratory
 *              Graduate School of Engineering Science, Osaka Univ., JAPAN
 *  Copyright (C) 2015,2016 by Embedded and Real-Time Systems Laboratory
 *              Graduate School of Information Science, Nagoya Univ., JAPAN
 * 
 *  上記著作権者は，以下の(1)～(4)の条件を満たす場合に限り，本ソフトウェ
 *  ア（本ソフトウェアを改変したものを含む．以下同じ）を使用・複製・改
 *  変・再配布（以下，利用と呼ぶ）することを無償で許諾する．
 *  (1) 本ソフトウェアをソースコードの形で利用する場合には，上記の著作
 *      権表示，この利用条件および下記の無保証規定が，そのままの形でソー
 *      スコード中に含まれていること．
 *  (2) 本ソフトウェアを，ライブラリ形式など，他のソフトウェア開発に使
 *      用できる形で再配布する場合には，再配布に伴うドキュメント（利用
 *      者マニュアルなど）に，上記の著作権表示，この利用条件および下記
 *      の無保証規定を掲載すること．
 *  (3) 本ソフトウェアを，機器に組み込むなど，他のソフトウェア開発に使
 *      用できない形で再配布する場合には，次のいずれかの条件を満たすこ
 *      と．
 *    (a) 再配布に伴うドキュメント（利用者マニュアルなど）に，上記の著
 *        作権表示，この利用条件および下記の無保証規定を掲載すること．
 *    (b) 再配布の形態を，別に定める方法によって，TOPPERSプロジェクトに
 *        報告すること．
 *  (4) 本ソフトウェアの利用により直接的または間接的に生じるいかなる損
 *      害からも，上記著作権者およびTOPPERSプロジェクトを免責すること．
 *      また，本ソフトウェアのユーザまたはエンドユーザからのいかなる理
 *      由に基づく請求からも，上記著作権者およびTOPPERSプロジェクトを
 *      免責すること．
 * 
 *  本ソフトウェアは，無保証で提供されているものである．上記著作権者お
 *  よびTOPPERSプロジェクトは，本ソフトウェアに関して，特定の使用目的
 *  に対する適合性も含めて，いかなる保証も行わない．また，本ソフトウェ
 *  アの利用により直接的または間接的に生じたいかなる損害に関しても，そ
 *  の責任を負わない．
 * 
 *  $Id$
 */

/*
 *		システムログタスクのコンポーネント記述ファイル
 */

/*
 *  システムログタスクのシグニチャ
 */
signature sLogTask {
	ER		flush([in] uint_t count);
};

/*
 *  システムログタスクの本体のセルタイプ
 */
[singleton]
celltype tLogTaskMain {
	entry	sTaskBody		eLogTaskBody;
	entry	sRoutineBody	eLogTaskTerminate;
	entry	sLogTask		eLogTask;

	call	sSerialPort		cSerialPort;	/* シリアルドライバとの接続 */
	call	snSerialPortManage	cnSerialPortManage;
											/* シリアルドライバ管理との接続 */
	call	sSysLog			cSysLog;		/* システムログ機能との接続 */
	call	sPutLog			cPutLog;		/* 低レベル出力との接続 */

	attr {
		RELTIM	interval;				/* システムログタスクの動作間隔 */
		RELTIM	flushWait;				/* フラッシュ待ちの単位時間 */
	};
};

/*
 *  システムログタスク（複合コンポーネント）のセルタイプ
 */
[singleton, active]
composite tLogTask {
	entry	sLogTask	eLogTask;		/* システムログタスク操作 */
	
	call	sSerialPort	cSerialPort;	/* シリアルドライバとの接続 */
	call	snSerialPortManage	cnSerialPortManage;
										/* シリアルドライバ管理との接続 */
	call	sSysLog		cSysLog;		/* システムログ機能との接続 */
	call	sPutLog		cPutLog;		/* 低レベル出力との接続 */

	attr {
		[omit] ATR		attribute = C_EXP("TA_ACT");	/* タスク属性 */
		[omit] PRI  	priority;		/* タスクの初期優先度 */
		[omit] size_t 	stackSize;		/* タスクのスタックサイズ */
		RELTIM		interval = 10000;	/* システムログタスクの動作間隔 */
		RELTIM		flushWait = 1000;	/* フラッシュ待ちの単位時間 */
	};

	cell tLogTaskMain LogTaskMain {
		/* 呼び口の結合 */
		cSerialPort        => composite.cSerialPort;
		cnSerialPortManage => composite.cnSerialPortManage;
		cSysLog            => composite.cSysLog;
		cPutLog            => composite.cPutLog;

		/* 属性の継承 */
		interval  = composite.interval;
		flushWait = composite.flushWait;
	};

	cell tTask Task {
		/* 呼び口の結合 */
		cTaskBody = LogTaskMain.eLogTaskBody;

		/* 属性の継承 */
		attribute = composite.attribute;
		priority  = composite.priority;
		stackSize = composite.stackSize;
	};

	cell tTerminateRoutine TerminateRoutine {
		/* 呼び口 */
		cTerminateRoutineBody = LogTaskMain.eLogTaskTerminate;
	};

	/* 受け口の結合 */
	composite.eLogTask => LogTaskMain.eLogTask;
};
