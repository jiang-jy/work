/*
 *		サンプルプログラム(1)のコンポーネント記述ファイル
 *
 *  $Id$
 */
/*
 *  カーネルオブジェクトの定義
 */
import(<kernel.cdl>);

/*
 *  ターゲット非依存のセルタイプの定義
 */
import("syssvc/tSerialPort.cdl");
import("syssvc/tSerialAdapter.cdl");
import("syssvc/tSysLog.cdl");
import("syssvc/tSysLogAdapter.cdl");
import("syssvc/tLogTask.cdl");
import("syssvc/tBanner.cdl");

/*
 *  ターゲット依存部の取り込み
 */
import("ntshell.cdl");
import_C("echonet.h");
/*
 *  「セルの組上げ記述」とは，"cell"で始まる行から，それに対応する"};"
 *  の行までのことを言う．
 */

/*
 *  システムログ機能の組上げ記述
 *
 *  システムログ機能を外す場合には，以下のセルの組上げ記述を削除し，コ
 *  ンパイルオプションに-DTOPPERS_OMIT_SYSLOGを追加すればよい．ただし，
 *  システムログタスクはシステムログ機能を使用するため，それも外すこと
 *  が必要である．また，システムログ機能のアダプタも外さなければならな
 *  い．tecsgenが警告メッセージを出すが，無視してよい．
 */
cell tSysLog SysLog {
	logBufferSize = 32;					/* ログバッファのサイズ */
	initLogMask = C_EXP("LOG_UPTO(LOG_NOTICE)");
										/* ログバッファに記録すべき重要度 */
	initLowMask = C_EXP("LOG_UPTO(LOG_EMERG)");
									   	/* 低レベル出力すべき重要度 */
	/* 低レベル出力との結合 */
	cPutLog = PutLogTarget.ePutLog;
};

/*
 *  C言語で記述されたアプリケーションから，TECSベースのシステムログ機能
 *  を呼び出すためのアダプタの組上げ記述
 *
 *  システムログ機能のサービスコール（syslog関数とsyslog_0関数～syslog_5
 *  関数以外のもの）ルをC言語で記述されたアプリケーションから呼び出さな
 *  い場合には，以下のセルの組上げ記述を削除すればよい．
 */
cell tSysLogAdapter SysLogAdapter {
	cSysLog = SysLog.eSysLog;
};

/*
 *  シリアルインタフェースドライバの組上げ記述
 *
 *  シリアルインタフェースドライバを外す場合には，以下のセルの組上げ記
 *  述を削除すればよい．ただし，システムログタスクはシリアルインタフェー
 *  スドライバを使用するため，それも外すことが必要である．また，シリア
 *  ルインタフェースドライバのアダプタも外さなければならない．
 */
cell tSerialPort SerialPort1 {
	receiveBufferSize = 256;			/* 受信バッファのサイズ */
	sendBufferSize    = 256;			/* 送信バッファのサイズ */

	/* ターゲット依存部との結合 */
	cSIOPort = SIOPortTarget1.eSIOPort;
	eiSIOCBR <= SIOPortTarget1.ciSIOCBR;	/* コールバック */
};

/*
 *  C言語で記述されたアプリケーションから，TECSベースのシリアルインタ
 *  フェースドライバを呼び出すためのアダプタの組上げ記述
 *
 *  シリアルインタフェースドライバのサービスコールをC言語で記述されたア
 *  プリケーションから呼び出さない場合には，以下のセルの組上げ記述を削
 *  除すればよい．
 */
cell tSerialAdapter SerialAdapter {
	cSerialPort[0] = SerialPort1.eSerialPort;
};

/*
 *  システムログタスクの組上げ記述
 *
 *  システムログタスクを外す場合には，以下のセルの組上げ記述を削除すれ
 *  ばよい．
 */
cell tLogTask LogTask {
	priority  = 3;					/* システムログタスクの優先度 */
	stackSize = LogTaskStackSize;	/* システムログタスクのスタックサイズ */

	/* シリアルインタフェースドライバとの結合 */
	cSerialPort        = SerialPort1.eSerialPort;
	cnSerialPortManage = SerialPort1.enSerialPortManage;

	/* システムログ機能との結合 */
	cSysLog = SysLog.eSysLog;

	/* 低レベル出力との結合 */
	cPutLog = PutLogTarget.ePutLog;
};

/*
 *  カーネル起動メッセージ出力の組上げ記述
 *
 *  カーネル起動メッセージの出力を外す場合には，以下のセルの組上げ記述
 *  を削除すればよい．
 */
cell tBanner Banner {
	/* 属性の設定 */
	targetName      = BannerTargetName;
	copyrightNotice = BannerCopyrightNotice;
};

//LightのTECS　CODE

/*
 * 
 *
 * 
 *
 *
 *　　　　　　　　　　　　　   　call Light　　　　    entry    call           entry
 *  +-------------+           +-------------+         +------------        +-------------+                     |------
 *  |             |           |             |         | tEchonet  |        |             |                     |
 *  |   tTask     | sTaskBody |   tTaskMain |sEchonet | Echonet   |slight  |  tLight     |                    |tLight
 *  |   Task      |-----------|>  TaskMain  |-------- |           |--------|>  Light     |              -------| Light
 *  |             |cTask      |             |         |           |        |             |(関数の定義)          |------
 *  |             |Body       |             |         |           |        |             |
 *  +-------------+           +-------------+         +------------       +-------------+                   other interface 
 *                        eTaskMain      cTaskMain            cEchonet     eLight
 *												                           light-echonet  interface 
 *						                              echonet interface                                       一般的照明用component interface						   	
 
//cfg file中的組件參數
 */                            

signature sEchonet{
	//ER main_initialize(void);
	
	void initialize(void);
	// ER main_get_timer(void);
	int getTimer(void);
	// ER main_progress([in]int interval);
	void progress([in] int interval);
	// ER main_recv_esv([in]T_EDATA *esv);
	//void ReciveService([in] const T_EDATA *esv, [in] int size);
	void ReciveService([in] const T_EDATA *esv);

	ER breakWait([in,size_is(len)] const uint8_t *brkdat,[in] int32_t len);
	//ER main_break_wait([in] const uint8_t *brkdat, [in] int32_t len);
	//ER main_timeout(void);
	void timeOut(void);
};

signature sLight{
	ER onOffPropertySet ([in] const uint8_t * src, [in]int size, [out]bool_t * anno);
	void OnPropertySet(void);
	void OffPropertySet(void);
 //echonet ``和light`的通信
// component 8-9以上. 
};

celltype tTaskMain{
	entry sTaskBody eTaskMain;
	call sEchonet cTaskMain;
};
cell tTaskMain TaskMain{
	cTaskMain = Echonet.eEchonet;
};

cell tTask Task{
	cTaskBody = TaskMain.eTaskMain;
	priority = 1;
	stackSize = 81920;
	attribute = C_EXP("TA_ACT");
};


celltype tEchonet{
	call sLight cEchonet;
	entry sEchonet eEchonet;
};

cell tEchonet Echonet{
	cEchonet = Light.eLight;
};


celltype tLight{
	entry sLight eLight;
	attr {
		
		uint8_t		eprpcd;			/* ECHONET Lite プロパティコード */
		//uint8_t   propertyCode;
		ATR			eprpatr;		/* ECHONET Lite プロパティ属性 */
		//uint8_t   propertyAttribute;
		uint8_t		eprpsz;			/* ECHONET Lite プロパティのサイズ */
		//uint8_t   propertySize;
		intptr_t	exinf;			/* ECHONET Lite プロパティの拡張情報 */
		//intptr_t	extendedInformation;	
		//EPRP_SETTER	*eprpset;		/* ECHONET Lite プロパティの設定関数 */
		//EPRP_GETTER	*eprpget;		/* ECHONET Lite プロパティの取得関数 */
		
		
	};
};
cell tLight Light{
		eprpcd=0;			/* ECHONET Lite プロパティコード */
		eprpatr=0;		 /*ECHONET Lite プロパティ属性 */
		eprpsz=0;			/* ECHONET Lite プロパティのサイズ */
		exinf=0;			/* ECHONET Lite プロパティの拡張情報 */
		//EPRP_SETTER	*eprpset;		/* ECHONET Lite プロパティの設定関数 */
		//EPRP_GETTER	*eprpget;		/* ECHONET Lite プロパティの取得関数 */
		
};
